`include "defines.vh"
module cpu_wrapper (
  input                   clock,
  input                   reset,
  input                   io_interrupt,
  input                   io_master_awready,
  output                  io_master_awvalid,
  output [`CPU_WIDTH-1:0] io_master_awaddr,
  output [           3:0] io_master_awid,
  output [           7:0] io_master_awlen,
  output [           2:0] io_master_awsize,
  output [           1:0] io_master_awburst,
  input                   io_master_wready,
  output                  io_master_wvalid,
  output [`CPU_WIDTH-1:0] io_master_wdata,
  output [           3:0] io_master_wstrb,
  output                  io_master_wlast,
  output                  io_master_bready,
  input                   io_master_bvalid,
  input  [           1:0] io_master_bresp,
  input  [           3:0] io_master_bid,
  input                   io_master_arready,
  output                  io_master_arvalid,
  output [`CPU_WIDTH-1:0] io_master_araddr,
  output [           3:0] io_master_arid,
  output [           7:0] io_master_arlen,
  output [           2:0] io_master_arsize,
  output [           1:0] io_master_arburst,
  output                  io_master_rready,
  input                   io_master_rvalid,
  input  [           1:0] io_master_rresp,
  input  [`CPU_WIDTH-1:0] io_master_rdata,
  input                   io_master_rlast,
  input  [           3:0] io_master_rid,
  output                  io_slave_awready,
  input                   io_slave_awvalid,
  input  [`CPU_WIDTH-1:0] io_slave_awaddr,
  input  [           3:0] io_slave_awid,
  input  [           7:0] io_slave_awlen,
  input  [           2:0] io_slave_awsize,
  input  [           1:0] io_slave_awburst,
  output                  io_slave_wready,
  input                   io_slave_wvalid,
  input  [`CPU_WIDTH-1:0] io_slave_wdata,
  input  [           3:0] io_slave_wstrb,
  input                   io_slave_wlast,
  input                   io_slave_bready,
  output                  io_slave_bvalid,
  output [           1:0] io_slave_bresp,
  output [           3:0] io_slave_bid,
  output                  io_slave_arready,
  input                   io_slave_arvalid,
  input  [`CPU_WIDTH-1:0] io_slave_araddr,
  input  [           3:0] io_slave_arid,
  input  [           7:0] io_slave_arlen,
  input  [           2:0] io_slave_arsize,
  input  [           1:0] io_slave_arburst,
  input                   io_slave_rready,
  output                  io_slave_rvalid,
  output [           1:0] io_slave_rresp,
  output [`CPU_WIDTH-1:0] io_slave_rdata,
  output                  io_slave_rlast,
  output [           3:0] io_slave_rid
);

  top u_top (
    .clock            (clock),
    .reset            (reset),
    .io_master_awready(io_master_awready),
    .io_master_awvalid(io_master_awvalid),
    .io_master_awaddr (io_master_awaddr),
    .io_master_awid   (io_master_awid),
    .io_master_awlen  (io_master_awlen),
    .io_master_awsize (io_master_awsize),
    .io_master_awburst(io_master_awburst),
    .io_master_wready (io_master_wready),
    .io_master_wvalid (io_master_wvalid),
    .io_master_wdata  (io_master_wdata),
    .io_master_wstrb  (io_master_wstrb),
    .io_master_wlast  (io_master_wlast),
    .io_master_bready (io_master_bready),
    .io_master_bvalid (io_master_bvalid),
    .io_master_bresp  (io_master_bresp),
    .io_master_bid    (io_master_bid),
    .io_master_arready(io_master_arready),
    .io_master_arvalid(io_master_arvalid),
    .io_master_araddr (io_master_araddr),
    .io_master_arid   (io_master_arid),
    .io_master_arlen  (io_master_arlen),
    .io_master_arsize (io_master_arsize),
    .io_master_arburst(io_master_arburst),
    .io_master_rready (io_master_rready),
    .io_master_rvalid (io_master_rvalid),
    .io_master_rresp  (io_master_rresp),
    .io_master_rdata  (io_master_rdata),
    .io_master_rlast  (io_master_rlast),
    .io_master_rid    (io_master_rid)
  );


endmodule
