module example();
    initial begin
        $display("Hello ysyx!");
    end
endmodule
